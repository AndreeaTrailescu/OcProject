library verilog;
use verilog.vl_types.all;
entity Iterator is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        i               : out    vl_logic_vector(3 downto 0)
    );
end Iterator;
